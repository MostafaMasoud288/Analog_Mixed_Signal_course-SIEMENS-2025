Simple RC Circuit

* Circuit Description

* Parameters
*** add line here ***
.PARAM CPAR=500p
* Signal sources
V1 1 0 PULSE(0V 1V 0 100n 100n 10u 20u)

* Circuit elements
R1 1 2 1k
C1 2 0 {CPAR}

* Initial conditions
.IC V(2)=0
* Analysis request
* Run transient for 40us with 100ns step
*** add line here ***
.TRAN 100n 40u
* Use parametric sweep for CPAR: 500p:500p:1.5n
*** add line here ***
*.STEP PARAM CPAR 500p 1.5n 500p
.STEP PARAM CPAR LIST 500p 1n 1.5n
* Measure rise time from 10% to 90%
.MEAS TRAN TRISE
+ TRIG when v(2) = 0.1 CROSS = 1
+ TARG WHEN V(2) = 0.9 CROSS = 1
*** add line here ***
.PRINT TRAN V(1) V(2)
.PLOT TRAN V(1) V(2)
*** add line here ***
.END
